
// REMOVE ME
