
`ifndef REGISTERS_SVH
`define REGISTERS_SVH


typedef struct packed {
    logic [23:0] Frequency;
    // feedback
    // amplitude
} OperatorConfiguration_t;


`endif
